module inv(a, y);
	input logic [0:0]a;
	output logic [0:0]y;	
	assign y = ~a;
endmodule 
